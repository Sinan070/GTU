library verilog;
use verilog.vl_types.all;
entity mips16 is
    port(
        clock           : in     vl_logic
    );
end mips16;
