library verilog;
use verilog.vl_types.all;
entity mips16Testbench is
end mips16Testbench;
