library verilog;
use verilog.vl_types.all;
entity cypher_detector_tb is
end cypher_detector_tb;
